netcdf udp_receive {
dimensions:
	dimS = 1 ;
	dimF = UNLIMITED ; // (12 currently)
variables:
	int index(dimF, dimS) ;
		index:units = "none" ;
		index:long_name = "received increment (from frame content)" ;
		index:frame_size_unit = "Byte" ;
		index:frame_size = 8192 ;
	int increment(dimF, dimS) ;
		increment:units = "none" ;
		increment:frame_size_unit = "Byte" ;
		increment:frame_size = 8192 ;

// global attributes:
		:library = "CImg_NetCDF" ;
		:library_version = "v0.8.4" ;
		:frame_size = 8192 ;
		:frame_size_unit = "BoF" ;
		:test_status = 0 ;
		:test_status_string = "fail" ;
		:mean_rate = 46.875f ;
		:mean_rate_unit = "MB/s" ;
		:elapsed_time = 2 ;
		:elapsed_time_unit = "ms" ;
		:expected_frame = 12 ;
		:expected_frame_unit = "frame" ;
		:received_frame = 12 ;
		:received_frame_unit = "frame" ;
		:total_drop = 2 ;
		:total_drop_unit = "drop" ;
		:total_index_drop = 107 ;
		:total_index_drop_unit = "index" ;
		:total_index_drop_percentage = 891.6667f ;
		:total_index_drop_percentage_unit = "%" ;
}

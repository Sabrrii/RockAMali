netcdf kernels
{
dimensions:

	kernel = 3; //UNLIMITED ;
	dimString=128;
variables:
	char kernel_name(kernel, dimString);
data:
	kernel_name = "0_discri", "1_discri_int2", "2_discri_int4";
}//kernels
netcdf udp_receive {
dimensions:
	dimS = 1 ;
	dimF = UNLIMITED ; // (121409 currently)
variables:
	int index(dimF, dimS) ;
		index:units = "none" ;
		index:long_name = "received index (from frame content)" ;
		index:frame_size_unit = "Byte" ;
		index:frame_size = 32768 ;
	int increment(dimF, dimS) ;
		increment:units = "none" ;
		increment:long_name = "received index (from frame content)" ;
		increment:frame_size_unit = "Byte" ;
		increment:frame_size = 32768 ;

// global attributes:
		:library = "CImg_NetCDF" ;
		:library_version = "v0.8.3" ;
		:frame_size = 32768 ;
		:frame_size_unit = "BoF" ;
		:test_status = 0 ;
		:test_status_string = "fail" ;
		:mean_rate = 77.49167f ;
		:mean_rate_unit = "MB/s" ;
		:elapsed_time = 49786 ;
		:elapsed_time_unit = "ms" ;
		:expected_frame = 123456 ;
		:expected_frame_unit = "frame" ;
		:received_frame = 121409 ;
		:received_frame_unit = "frame" ;
		:total_drop = 134 ;
		:total_drop_unit = "drop" ;
		:total_index_drop = 2048 ;
		:total_index_drop_unit = "index" ;
		:total_index_drop_percentage = 1.658891f ;
		:total_index_drop_percentage_unit = "%" ;
}

netcdf result_sequential {
dimensions:
	dimS = 8192 ;
	dimF = UNLIMITED ; // (23 currently)
variables:
	int signal(dimF, dimS) ;
		signal:units = "digit" ;
		signal:long_name = "GPU discri signal" ;
		signal:kernel = "CDataProcessorGPU_discri_opencl_int4" ;

// global attributes:
		:kernel = "CDataProcessorGPU_discri_opencl_int4" ;
}

netcdf result_sequential {
dimensions:
	dimS = 1 ;
	dimF = UNLIMITED ; // (23 currently)
variables:
	int E(dimF, dimS) ;
		E:units = "digit" ;
		E:long_name = "energy" ;
		E:kernel = "CDataProcessorGPU_discri_opencl_int4" ;

// global attributes:
		:kernel = "CDataProcessorGPU_discri_opencl_int4" ;
}

netcdf RockAMali.parameters {//written in NetCDF CDL language
  :institution = "GANIL";
  :title = "RockAMali parameters";
  :comment = "source of parameters for RockAMali processing program";
  :history = "";
  :version = "v0.0.1";

dimensions:
//  dim_string=64;
//  dim_=unlimited;

//variable declaration and attributes
variables:
//signal
  int signal;
     signal:long_name="signal graph (activated if >0)";
     signal:nb_tB_long_name="baseline time";
     signal:nb_tB= 1234; 
     signal:nb_tA_long_name="peak time"; 
     signal:nb_tA= 10; 
     signal:tau_long_name="time decrease";
     signal:tau= 500;
     signal:A_long_name="Amplitude";
     signal:A= 2345;
     signal:B_long_name="Baseline";
     signal:B= 23;
//Generator Random
     signal:rand_min=0;
     signal:rand_max=65535;
//Generator full_random
     signal:noise=0.2;//12.3;
//! \todo noise_ampl instead of min_Amp and max_Amp, same for tau, tA, tB (+B)
     signal:min_tB=1234;
     signal:max_tB=1235;
     signal:noise_tA_long_name="peak noise time amplitude"; 
     signal:noise_tA=2;
     signal:noise_B=3;
     signal:noise_A=12;
     signal:min_tau=500;
     signal:max_tau=501;


//trapezoid filter
  int trapezoid;
    trapezoid:long_name="trapezoid filter (activated if >0)";
    trapezoid:k_long_name= "increase size";
    trapezoid:k= 200;
    trapezoid:k_units= "pixel";
    trapezoid:m_long_name= "plateau size";
    trapezoid:m= 50;
    trapezoid:m_units= "pixel";
    trapezoid:alpha_long_name= "";
    trapezoid:alpha= 0.99800199866733306675;
    trapezoid:alpha_units= "";
    trapezoid:n= 34;
    trapezoid:q= 211;
    trapezoid:q_long_name= "Q computing delay";
    trapezoid:threshold=3.4;
    trapezoid:fraction=0.2;
    trapezoid:Tm=20;

//data value
data:
//signal
  signal=1;
//trapezoid filter
  trapezoid=1;
}


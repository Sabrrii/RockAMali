netcdf profiling_process {
dimensions:
	dim1 = 1 ;
	dimF = UNLIMITED ; // (23 currently)
variables:
	int iteration(dimF, dim1) ;
		iteration:units = "us" ;
		iteration:kernel = "CDataProcessor_Max_Min" ;
		iteration:frame_size = 8192 ;
	int storage(dimF, dim1) ;
		storage:units = "us" ;
		storage:storage = "CDataStore" ;
		storage:frame_size = 8192 ;
	int process_sequential_elapsed_time ;
		process_sequential_elapsed_time:units = "us" ;
		process_sequential_elapsed_time:profiling = "CProfilingSequential" ;
	int process_sequential_elapsed_time_per_iteration ;
		process_sequential_elapsed_time_per_iteration:units = "us" ;
		process_sequential_elapsed_time_per_iteration:profiling = "CProfilingSequential" ;

// global attributes:
		:process_sequential = "v0.7.3r" ;
		:CImg_NetCDF = "v0.8.3" ;
		:CParameterNetCDF = "v0.5.0" ;
		:NcTypeInfo = "v0.1.4" ;
		:kernel = "CDataProcessor_Max_Min" ;
		:profiling = "CProfilingSequential" ;
		:process_sequential_elapsed_time = 23017 ;
		:process_sequential_elapsed_time_units = "us" ;
		:process_sequential_elapsed_time_per_iteration = 1000 ;
}

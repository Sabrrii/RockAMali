netcdf pac_signal_parameters {
dimensions:
	dim1 = 1 ;
	dimF = UNLIMITED ; // (23 currently)
variables:
	int A(dimF, dim1) ;
		A:units = "digit" ;
		A:long_name = "amplitude" ;
		A:generator_ = "CDataGenerator_Peak" ;
		A:generator = "CDataGenerator_Full_Random" ;
	int B(dimF, dim1) ;
		B:units = "digit" ;
		B:long_name = "baseline" ;
		B:generator_ = "CDataGenerator_Peak" ;
		B:generator = "CDataGenerator_Full_Random" ;
	int tB(dimF, dim1) ;
		tB:units = "tic (10ns)" ;
		tB:long_name = "baseline duration" ;
		tB:generator_ = "CDataGenerator_Peak" ;
		tB:generator = "CDataGenerator_Full_Random" ;
	int tA(dimF, dim1) ;
		tA:units = "tic (10ns)" ;
		tA:long_name = "increase duration" ;
		tA:generator_ = "CDataGenerator_Peak" ;
		tA:generator = "CDataGenerator_Full_Random" ;
	int Tau(dimF, dim1) ;
		Tau:units = "tic (10ns)" ;
		Tau:long_name = "exponential decrease" ;
		Tau:generator_ = "CDataGenerator_Peak" ;
		Tau:generator = "CDataGenerator_Full_Random" ;
	int E(dimF, dim1) ;
		E:units = "digit" ;
		E:long_name = "energy (computed using E=A-B)" ;
		E:generator_ = "CDataGenerator_Peak" ;
		E:generator = "CDataGenerator_Full_Random" ;

// global attributes:
		:architecture = "x86_64" ;
		:signal_noise_min = -0.1f ;
		:signal_noise_max = 0.1f ;
}

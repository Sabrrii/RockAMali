netcdf profiling_gpu {
dimensions:
	dimP = 1 ;
	dimF = UNLIMITED ; // (23 currently)
variables:
	int kernel_elapsed_time(dimF, dimP) ;
		kernel_elapsed_time:units = "us" ;
		kernel_elapsed_time:kernel = "CDataProcessorGPU_discri_opencl_int4" ;

// global attributes:
		:architecture = "ARM64" ;
}

netcdf udp_receive {
dimensions:
	dimS = 1 ;
	dimF = UNLIMITED ; // (12289 currently)
variables:
	int index(dimF, dimS) ;
		index:units = "none" ;
		index:long_name = "received index (from frame content)" ;
		index:frame_size_unit = "Byte" ;
		index:frame_size = 32768 ;

// global attributes:
		:library = "CImg_NetCDF" ;
		:library_version = "v0.8.3" ;
		:frame_size = 32768 ;
		:frame_size_unit = "BoF" ;
		:test_status = 0 ;
		:test_status_string = "fail" ;
		:mean_rate = 38.66319f ;
		:mean_rate_unit = "MB/s" ;
		:elapsed_time = 9978 ;
		:elapsed_time_unit = "ms" ;
		:expected_frame = 12345 ;
		:expected_frame_unit = "frame" ;
		:received_frame = 12289 ;
		:received_frame_unit = "frame" ;
		:total_drop = 21 ;
		:total_drop_unit = "drop" ;
		:total_index_drop = 57 ;
		:total_index_drop_unit = "index" ;
		:total_index_drop_percentage = 0.4617254f ;
		:total_index_drop_percentage_unit = "%" ;
}
